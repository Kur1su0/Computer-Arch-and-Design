CAD_lib.lab9_register_decoder(behav) :5:
CAD_lib.lab9_regReadWrite(mixed) :32:
