CAD_lib.reg(mixed) :32:
