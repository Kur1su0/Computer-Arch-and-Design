--
-- VHDL Architecture CAD_lib.lab3_fetch_unit.behav
--
-- Created:
--          by - W.UNKNOWN (DESKTOP-86TQKQ1)
--          at - 22:55:02 02/22/2021
--
-- using Mentor Graphics HDL Designer(TM) 2018.2 (Build 19)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY lab3_fetch_unit IS
END ENTITY lab3_fetch_unit;

--
ARCHITECTURE behav OF lab3_fetch_unit IS
BEGIN
END ARCHITECTURE behav;

