CAD_lib.reg(mixed) :32:
CAD_lib.reg(mixed) :5:
CAD_lib.func_reg(behav) rtlc_no_parameters
