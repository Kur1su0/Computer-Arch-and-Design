CAD_lib.mux_2_to_1(mixed) :32:
