--
-- VHDL Architecture CAD_lib.inc.mixed
--
-- Created:
--          by - W.UNKNOWN (DESKTOP-86TQKQ1)
--          at - 20:34:13 02/12/2021
--
-- using Mentor Graphics HDL Designer(TM) 2018.2 (Build 19)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY inc IS
END ENTITY inc;

--
ARCHITECTURE mixed OF inc IS
BEGIN
END ARCHITECTURE mixed;

