CAD_lib.reg(mixed) :32:
CAD_lib.reg(mixed) :5:
CAD_lib.func_reg(behav) rtlc_no_parameters
CAD_lib.lab9_register_decoder(behav) :5:
CAD_lib.lab9_regReadWrite(mixed) :32:
