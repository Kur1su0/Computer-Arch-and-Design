--
-- VHDL Architecture CAD_lib.lab8_writeback.mixed
--
-- Created:
--          by - W.UNKNOWN (DESKTOP-86TQKQ1)
--          at - 02:53:40 04/ 4/2021
--
-- using Mentor Graphics HDL Designer(TM) 2018.2 (Build 19)
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY lab8_writeback IS
END ENTITY lab8_writeback;

--
ARCHITECTURE mixed OF lab8_writeback IS
BEGIN
END ARCHITECTURE mixed;

