CAD_lib.lab9_register_decoder(behav) :5:
